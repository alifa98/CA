--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   00:03:40 12/24/2019
-- Design Name:   
-- Module Name:   C:/Users/aliwin/Desktop/VHDL/Memory/CAM_TB.vhd
-- Project Name:  Memory
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: CAM
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY CAM_TB IS
END CAM_TB;
 
ARCHITECTURE behavior OF CAM_TB IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT CAM
    PORT(
         clock : IN  std_logic;
         rw : IN  std_logic;
         reset : IN  std_logic;
         data : IN  std_logic_vector(2 downto 0);
         match : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clock : std_logic := '0';
   signal rw : std_logic := '0';
   signal reset : std_logic := '0';
   signal data : std_logic_vector(2 downto 0) := (others => '0');

 	--Outputs
   signal match : std_logic;

   -- Clock period definitions
   constant clock_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: CAM PORT MAP (
          clock => clock,
          rw => rw,
          reset => reset,
          data => data,
          match => match
        );

   -- Clock process definitions
   clock_process :process
   begin
		clock <= '0';
		wait for clock_period/2;
		clock <= '1';
		wait for clock_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 105 ns;	

      wait for clock_period*10;
		reset <= '1';
		rw <= '1';
		data <= "101";

      wait for clock_period*10;
		rw <= '0';
		data <= "111";

      wait for clock_period*10;
		rw <= '0';
		data <= "101";

      wait for clock_period*10;
		rw <= '1';
		data <= "111";

      wait for clock_period*10;
		rw <= '0';
		data <= "111";

      wait for clock_period*10;
		reset <= '0';
		rw <= '1';
		data <= "101";

      wait for clock_period*10;
		reset <= '1';
		rw <= '0';
		data <= "101";

      wait for clock_period*10;
		rw <= '1';
		data <= "001";   

		wait for clock_period*10;
		rw <= '0';
		data <= "001";
		
		
      wait;
   end process;

END;

